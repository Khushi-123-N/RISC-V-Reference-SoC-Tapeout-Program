﻿	imescale 1ns/1ps

module example_module_tb;

reg clk;
reg rst;
reg [3:0] in_data;
wire [3:0] out_data;

example_module uut (
    .clk(clk),
    .rst(rst),
    .in_data(in_data),
    .out_data(out_data)
);

initial begin
    clk = 0;
    forever #5 clk = ~clk; // 100MHz clock
end

initial begin
    rst = 1;
    in_data = 4'b0000;
    #10;
    rst = 0;
    #10;
    in_data = 4'b1010;
    #20;
    in_data = 4'b0101;
    #20;
    ;
end

endmodule
